`ifndef AHBRAM_TESTS_SV
`define AHBRAM_TSETS_SV

`include "ahbram_base_test.sv"
`include "ahbram_smoke_test.sv"
`include "ahbram_diff_hsize_test.sv"
`include "ahbram_diff_haddr_test.sv"
`include "ahbram_reset_w2r_test.sv"
`include "ahbram_haddr_word_unaligned_test.sv"
`include "ahbram_htrans_test.sv"
 

`endif 