`ifndef AHB_PKG_SV
`define AHB_PKG_SV

package ahb_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "ahb_defines.svh"
    `include "ahb_types.sv"
    `include "ahb_configuration.sv" 
    `include "ahb_agent_configuration.sv"
    `include "ahb_transaction.sv"  
    `include "ahb_sequencer.sv"  
    `include "ahb_driver.sv"  
    `include "ahb_monitor.sv"  
    `include "ahb_master_transaction.sv"  
    `include "ahb_master_driver.sv"  
    `include "ahb_master_monitor.sv"  
    `include "ahb_master_sequencer.sv"  
    `include "ahb_master_agent.sv"  
    `include "ahb_sequence_lib.svh"

endpackage


`endif 
