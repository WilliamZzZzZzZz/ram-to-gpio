`ifndef RKV_GPIO_SEQ_LIB_SVH
`define RKV_GPIO_SEQ_LIB_SVH

`include "rkv_gpio_element_sequences.svh"
`include "rkv_gpio_base_virtual_sequence.sv"
`include "rkv_gpio_portout_set_virt_seq.sv"
`include "rkv_gpio_interrupt_virt_seq.sv"
`include "rkv_gpio_masked_virt_seq.sv"


`endif
