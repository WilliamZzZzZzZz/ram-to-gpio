`ifndef AHB_SEQUENCE_LIB_SV
`define AHB_SEQUENCE_LIB_SV

`include "ahb_base_sequence.sv"
`include "ahb_master_single_sequence.sv"

`endif 