`ifndef RKV_GPIO_TESTS_SVH
`define RKV_GPIO_TESTS_SVH

`include "rkv_gpio_base_test.sv"
`include "rkv_gpio_portout_set_test.sv"
`include "rkv_gpio_interrupt_test.sv"
`include "rkv_gpio_masked_test.sv"
`include "rkv_gpio_output_enable_test.sv"

`endif // RKV_GPIO_TESTS_SVH
